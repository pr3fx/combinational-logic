module full_adder (
                   input logic  a, b,
                   output logic s, cout
                   );
   

endmodule // full_adder
