module mux4 (
             input logic [3:0] a,
             output logic      y
             );
   
endmodule // mux4
