module cla
  #(parameter width=16)
   (input logic              cin,
    input logic [width-1:0]  a, b,
    output logic [width-1:0] s,
    output logic             cout);

endmodule // cla
