module prefix_adder
  #(parameter width=8)
   (input logic              cin,
    input logic [width-1:0]  a, b,
    output logic             cout,
    output logic [width-1:0] s);

endmodule // prefix_adder
